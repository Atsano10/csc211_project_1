`timescale 1ns/1ps

module tb_toUpper;

reg [7:0] a;
wire [7:0] b;

toUpper dut (.a(a), .b(b));

initial begin
    $dumpfile("toUpper.vcd");
    $dumpvars(0, tb_toUpper);
    
    // (
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b00101000; #26;
    // H
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01001000; #26;
    // .
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b10110111; #26;
    // f
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b10000011; #26;
    // |
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01111100; #26;
    // DC4
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b00010100; #26;
    // ë
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b11101011; #26;
    // a
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01100001; #26;
    // A
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01000001; #26;
    // z
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01111010; #26;
    // G
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01000111; #26;
    // m
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01101101; #26;
    // '
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b10010010; #26;
    // 0
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b00110000; #26;
    // Ï
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b11001111; #26;
    // : 
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b00111010; #26;
    // {
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01111011; #26;
    // ”
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b10010100; #26;
    // DEL
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01111111; #26;

    #50 $finish;
end

endmodule
