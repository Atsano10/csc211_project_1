module tb_toUpper;

reg [7:0] a;
wire [7:0] b;

toUpper dut (.a(a), .b(b));

initial begin
    $dumpfile("toUpper.vcd");
    $dumpvars(0, tb_toUpper);
    
    // (
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b00101000; #15;
    // H
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01001000; #15;
    // .
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b10110111; #15;
    // f
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b10000011; #15;
    // |
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01111100; #15;
    // DC4
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b00010100; #15;
    // ë
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b11101011; #15;
    // a
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01100001; #15;
    // A
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01000001; #15;
    // z
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01111010; #15;
    // G
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01000111; #15;
    // m
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01101101; #15;
    // '
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b10010010; #15;
    // 0
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b00110000; #15;
    // Ï
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b11001111; #15;
    // : 
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b00111010; #15;
    // {
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01111011; #15;
    // ”
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b10010100; #15;
    // DEL
    {a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]} = 8'b01111111; #15;

    #50 $finish;
end

endmodule